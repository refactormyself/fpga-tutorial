`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
//////////////////////////////////////////////////////////////////////////////////


module AndCircuit(
    output out,
    input in1,
    input in2
    );
    
    and(out, in1, in2);
endmodule
