`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//This gives as output the 1's compliment of the input 
// Does a compliment of all the bits
//////////////////////////////////////////////////////////////////////////////////


module OnesCompliment(
    input [7:0] In,
    output [7:0] Out
    );
    assign Out = ~In;
endmodule
