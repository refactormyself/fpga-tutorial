`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
//////////////////////////////////////////////////////////////////////////////////


module MyAndGate(
    input In1,
    input In2,
    input Out
    );
    
    assign Out = In1 & In2;
endmodule
