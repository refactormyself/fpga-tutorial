`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
//////////////////////////////////////////////////////////////////////////////////


module MyFullAdder(
     input  A,
     input  B,
     input  Cin,
     output S,
     output Cout
     );
     assign S = A^B^Cin;
     assign Cout = (A&B) | (A&Cin) | (B&Cin);
endmodule
