`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
//////////////////////////////////////////////////////////////////////////////////


module AndOrCircuit(
    output out,
    input in1,
    input in2,
    input in3
    );
    
    wire andOut;
    and(andOut, in1, in2);
    or(out, in3, andOut);
endmodule
